    Mac OS X            	   2  
     <                                      ATTR      <   �   t                  �   .  %com.apple.metadata:kMDItemWhereFroms    �   F  com.apple.quarantine bplist00�P                            q/0001;5a2019a2;Google\x20Chrome;15B73808-DB68-4F82-80F8-6C1D0AEF9D51 