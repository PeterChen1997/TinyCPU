    Mac OS X            	   2  
     <                                      ATTR      <   �   t                  �   .  %com.apple.metadata:kMDItemWhereFroms    �   F  com.apple.quarantine bplist00�P                            q/0001;5a201994;Google\x20Chrome;E42FA135-7769-4772-A3C7-925C4355E28A 