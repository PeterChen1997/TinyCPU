    Mac OS X            	   2  
     <                                      ATTR      <   �   t                  �   .  %com.apple.metadata:kMDItemWhereFroms    �   F  com.apple.quarantine bplist00�P                            q/0001;5a2019d4;Google\x20Chrome;74DBC9EA-3E4E-49D2-841F-55647A896712 