    Mac OS X            	   2  
     <                                      ATTR      <   �   t                  �   .  %com.apple.metadata:kMDItemWhereFroms    �   F  com.apple.quarantine bplist00�P                            q/0001;5a2019d2;Google\x20Chrome;EEF700D7-72EF-4C39-8D9E-514E1917163F 