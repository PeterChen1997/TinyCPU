    Mac OS X            	   2  
     <                                      ATTR      <   �   t                  �   .  %com.apple.metadata:kMDItemWhereFroms    �   F  com.apple.quarantine bplist00�P                            q/0001;5a20198f;Google\x20Chrome;E23CE587-E780-4B19-AB13-188446B71734 