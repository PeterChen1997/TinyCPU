    Mac OS X            	   2  
     <                                      ATTR      <   �   t                  �   .  %com.apple.metadata:kMDItemWhereFroms    �   F  com.apple.quarantine bplist00�P                            q/0001;5a2019c3;Google\x20Chrome;49D7B0CC-55AD-46BC-B1DF-D170E8939F92 