    Mac OS X            	   2  
     <                                      ATTR      <   �   t                  �   .  %com.apple.metadata:kMDItemWhereFroms    �   F  com.apple.quarantine bplist00�P                            q/0001;5a201976;Google\x20Chrome;E771EA7C-42C3-41C3-B4E3-90BBFE5ED8FF 