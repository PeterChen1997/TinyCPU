    Mac OS X            	   2  
     <                                      ATTR      <   �   t                  �   .  %com.apple.metadata:kMDItemWhereFroms    �   F  com.apple.quarantine bplist00�P                            q/0001;5a201981;Google\x20Chrome;9AD9745E-B3F2-4B16-86A6-E4B7A284BC2C 