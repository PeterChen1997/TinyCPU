    Mac OS X            	   2  
     <                                      ATTR      <   �   t                  �   .  %com.apple.metadata:kMDItemWhereFroms    �   F  com.apple.quarantine bplist00�P                            q/0001;5a2019af;Google\x20Chrome;996861FE-5FDF-4B74-87F2-09FBA790C694 