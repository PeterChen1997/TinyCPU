    Mac OS X            	   2  
     <                                      ATTR      <   �   t                  �   .  %com.apple.metadata:kMDItemWhereFroms    �   F  com.apple.quarantine bplist00�P                            q/0001;5a2019bb;Google\x20Chrome;3C915FFA-26D5-458B-80C3-A42CB7C112EE 